library	ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity s_dcd is
	port(nr:in std_logic_vector(8 downto 0);
	x3,x2,x1,x0:out std_logic_vector(6 downto 0));
end s_dcd;
architecture f1 of s_dcd is
begin	   
	
	process(nr)
	variable dec:std_logic_vector(6 downto 0);
	begin
		case nr is
			when "000000000"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0000001";--0
			when "000000001"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="1001111";--1
			when "000000010"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0010010";--2
			when "000000011"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0000110";--3 
			when "000000100"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="1001100";--4	
			when "000000101"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0100100";--5
			when "000000110"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0100000";--6
			when "000000111"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0001111";--7
			when "000001000"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0000000";--8
			when "000001001"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0001000";--9
			when "000001010"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0000001"; --10
			when "000001011"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="1001111"; --11
			when "000001100"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="1101101"; --12
			when "000001101"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0000110";--13
			when "000001110"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="1001100";--14
			when "000001111"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0100100";--15
			when "000010000"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0100000";--16  
			when "000010001"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0001111";--17
			when "000010010"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0000000";--18
			when "000010011"=>x3<="0000001";x2<="0000001";x1<="1001111";x0<="0001000";--19
			when "000010100"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0000001";--20
			when "000010101"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="1001111";--21
			when "000010110"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0010010";--22
			when "000010111"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0000110";--23
			when "000011000"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="1001100";--24
			when "000011001"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0100100";--25
			when "000011010"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0100000";--26
			when "000011011"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0001111";--27
			when "000011100"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0000000";--28
			when "000011101"=>x3<="0000001";x2<="0000001";x1<="0010010";x0<="0001000";--29  
			when "000011110"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0000001";--30
			when "000011111"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="1001111";--31
			when "000100000"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0010010";--32
			when "000100001"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0000110";--33
			when "000100010"=>x3<="0000001";x2<="0000001";x1<="1001100";x0<="1001100";--34
			when "000100011"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0100100";--35																				 --35
		    when "000100100"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0100000";--36
			when "000100101"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0001111";--37
		    when "000100110"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0000000";--38
			when "000100111"=>x3<="0000001";x2<="0000001";x1<="0000110";x0<="0001000";--39
			when "000101000"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0000001";--40
			when "000101001"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="1001111";--41
			when "000101010"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0010010";--42	 
			when "000101011"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0000110";--43
			when "000101100"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="1001100";--44
			when "000101101"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0100100";--45
			when "000101110"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0100000";--46
			when "000101111"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0001111";--47
			when "000110000"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0000000";--48
			when "000110001"=>x3<="0000001";x2<="0000001";x1<="0001100";x0<="0001000";--49
			when "000110010"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0000001";--50  
			when "000110011"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="1001111";--51
			when "000110100"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0010010";--52
			when "000110101"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0000110";--53
			when "000110110"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="1001100";--54
			when "000110111"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0100100";--55
			when "000111000"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0100000";--56
			when "000111001"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0001111";--57
			when "000111010"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0000000";--58
			when "000111011"=>x3<="0000001";x2<="0000001";x1<="0100100";x0<="0001000";--59
			when "000111100"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0000001";--60
			when "000111101"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="1001111";--61
			when "000111110"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0010010";--62
			when "000111111"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0000110";--63
			when "001000000"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="1001100";--64
			when "001000001"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0100100";--65
			when "001000010"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0100000";--66
			when "001000011"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0001111";--67
			when "001000100"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0000000";--68
			when "001000101"=>x3<="0000001";x2<="0000001";x1<="0100000";x0<="0001000";--69 
			when "001000110"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0000001";--70
			when "001000111"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="1001111";--71
			when "001001000"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0010010";--72
			when "001001001"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0000110";--73
			when "001001010"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="1001100";--74
			when "001001011"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0100100";--75
			when "001001100"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0100000";--76
			when "001001101"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0001111";--77
			when "001001110"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0000000";--78
			when "001001111"=>x3<="0000001";x2<="0000001";x1<="0001111";x0<="0001000";--79
			when "001010000"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0000001";--80
			when "001010001"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="1001111";--81
			when "001010010"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0010010";--82
			when "001010011"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0000110";--83
			when "001010100"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="1001100";--84
			when "001010101"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0100100";--85
			when "001010110"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0100000";--86
			when "001010111"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0001111";--87
			when "001011000"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0000000";--88
			when "001011001"=>x3<="0000001";x2<="0000001";x1<="0000000";x0<="0001000";--89 
			when "001011010"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0000001";--90
			when "001011011"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="1001111";--91
			when "001011100"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0010010";--92
			when "001011101"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0000110";--93
			when "001011110"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="1001100";--94
			when "001011111"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0100100";--95
			when "001100000"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0100000";--96
			when "001100001"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0001111";--97
			when "001100010"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0000000";--98
			when "001100011"=>x3<="0000001";x2<="0000001";x1<="0001000";x0<="0001000";--99
			when "001100100"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0000001";--100
			when "001100101"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="1001111";--101
			when "001100110"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0010010";--102
			when "001100111"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0000110";--103
			when "001101000"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="1001100";--104
			when "001101001"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0100100";--105
			when "001101010"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0100000";--106
			when "001101011"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0001111";--107
			when "001101100"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0000000";--108
			when "001101101"=>x3<="0000001";x2<="1001111";x1<="0000001";x0<="0001000";--109
			when "001101110"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0000001";--110
			when "001101111"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0000001";--111
			when "001110000"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0010010";--112
			when "001110001"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0000110";--113
			when "001110010"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="1001100";--114
			when "001110011"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0100100";--115
			when "001110100"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0100000";--116
			when "001110101"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0001111";--117
			when "001110110"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0000000";--118
			when "001110111"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0001000";--119
			when "001111000"=>x3<="0000001";x2<="1001111";x1<="1001111";x0<="0000001";--120
			when "001111001"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="0000001";--121
			when "001111010"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="0010010";--122
			when "001111011"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="0000110";--123
			when "001111100"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="1001100";--124
			when "001111101"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="0100100";--125
			when "001111110"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="0100000";--126
			when "001111111"=>x3<="0000001";x2<="1001111";x1<="0010010";x0<="0001111";--127
			
			when "010000000"=>x3<="0000001";x2<="0000001";x1<="0000001";x0<="0000001";--0	
			when "010000001"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="0001111";-- -127
			when "010000010"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="0100000";-- -126
			when "010000011"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="0100100";-- -125
			when "010000100"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="1001100";-- -124 
			when "010000101"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="0000110";--  -123
			when "010000110"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="0010010";--  -122
			when "010000111"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="1001111";--  -121
			when "010001000"=>x3<="1111110";x2<="1001111";x1<="0010010";x0<="0000001";--  -120
			when "010001001"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0001000";--  -119
			when "010001010"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0000000";--  -118
			when "010001011"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0001111";--  -117
			when "010001100"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0100000";--  -116
			when "010001101"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0100100";--  -115
			when "010001110"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="1001100";--  -114
			when "010001111"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0000110";--  -113
			when "010010000"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0010010";--  -112  
			when "010010001"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="1001111";--  -111
			when "010010010"=>x3<="1111110";x2<="1001111";x1<="1001111";x0<="0000001";--  -110
			when "010010011"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0001000";--  -109
			when "010010100"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0000000";--  -108
			when "010010101"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0001111";--	 -107
			when "010010110"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0100000";--  -106
			when "010010111"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0100100";--  -105
			when "010011000"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="1001100";--  -104
			when "010011001"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0000110";--  -103
			when "010011010"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0010010";--  -102
			when "010011011"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="1001111";--  -101
			when "010011100"=>x3<="1111110";x2<="1001111";x1<="0000001";x0<="0000001";--  -100
			when "010011101"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0001000";--  -99  
			when "010011110"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0000000";--  -98
			when "010011111"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0001111";--  -97
			when "010100000"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0100000";--  -96
			when "010100001"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0100100";--  -95
			when "010100010"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="1001100";--  -94
			when "010100011"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0000110";--  -93																				 --35
		    when "010100100"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0010010";--  -92
			when "010100101"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="1001111";--  -91
		    when "010100110"=>x3<="1111110";x2<="0000001";x1<="0000100";x0<="0000001";--  -90
			when "010100111"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0001000";--  -89
			when "010101000"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0000000";--  -88
			when "010101001"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0001111";--  -87
			when "010101010"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0100000";--  -86 
			when "010101011"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0100100";--  -85
			when "010101100"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="1001100";--  -84
			when "010101101"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0000110";--  -83
			when "010101110"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0010010";--  -82
			when "010101111"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="1001111";--  -81
			when "010110000"=>x3<="1111110";x2<="0000001";x1<="0000000";x0<="0000001";--  -80
			when "010110001"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0001000";--  -79
			when "010110010"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0000000";--  -78
			when "010110011"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0001111";--  -77
			when "010110100"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0100000";--  -76
			when "010110101"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0100100";--  -75
			when "010110110"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="1001100";--  -74
			when "010110111"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0000110";--  -73
			when "010111000"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0010010";--  -72
			when "010111001"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="1001111";--  -71
			when "010111010"=>x3<="1111110";x2<="0000001";x1<="0001111";x0<="0000001";--  -70
			when "010111011"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0001000";--  -69
			when "010111100"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0000000";--  -68
			when "010111101"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0001111";--  -67
			when "010111110"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0100000";--  -66
			when "010111111"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0100100";--  -65
			when "011000000"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="1001100";--  -64
			when "011000001"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0000110";--  -63
			when "011000010"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0010010";--  -62
			when "011000011"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="1001111";--  -61
			when "011000100"=>x3<="1111110";x2<="0000001";x1<="0100000";x0<="0000001";--  -60
			when "011000101"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0001000";--  -59 
			when "011000110"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0000000";--  -58
			when "011000111"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="1110000";--  -57
			when "011001000"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0100000";--  -56
			when "011001001"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0100100";--  -55
			when "011001010"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="1001100";--  -54
			when "011001011"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0000110";--  -53
			when "011001100"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0010010";--  -52
			when "011001101"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="1001111";--  -51
			when "011001110"=>x3<="1111110";x2<="0000001";x1<="0100100";x0<="0000001";--  -50
			when "011001111"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0001000";--  -49
			when "011010000"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0000000";--  -48
			when "011010001"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="1110000";--  -47
			when "011010010"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0100000";--  -46
			when "011010011"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0100100";--  -45
			when "011010100"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="1001100";--  -44
			when "011010101"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0000110";--  -43
			when "011010110"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0010010";--  -42
			when "011010111"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="1001111";--  -41
			when "011011000"=>x3<="1111110";x2<="0000001";x1<="1001100";x0<="0000001";--  -40
			when "011011001"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0001000";--  -39 
			when "011011010"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0000000";--  -38
			when "011011011"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0001111";--  -37
			when "011011100"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0100000";--  -36
			when "011011101"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0100100";--  -35
			when "011011110"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="1001100";--  -34
			when "011011111"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0000110";--  -33
			when "011100000"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0100010";--  -32
			when "011100001"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="1001111";--  -31 
			when "011100010"=>x3<="1111110";x2<="0000001";x1<="0000110";x0<="0000001";--  -30
			when "011100011"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0001000";--  -29
			when "011100100"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0000000";--  -28
			when "011100101"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0001111";--  -27
			when "011100110"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0100000";--  -26
			when "011100111"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0100100";--  -25
			when "011101000"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="1001100";--  -24
			when "011101001"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0000110";--  -23
			when "011101010"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0010010";--  -22
			when "011101011"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="1001111";--  -21
			when "011101100"=>x3<="1111110";x2<="0000001";x1<="0010010";x0<="0000001";--  -20
			when "011101101"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0001000";--  -19
			when "011101110"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0000000";--  -18
			when "011101111"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0001111";--  -17
			when "011110000"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0100000";--  -16
			when "011110001"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0100100";--  -15
			when "011110010"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="1001100";--  -14
			when "011110011"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0000110";--  -13
			when "011110100"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0010010";--  -12
			when "011110101"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="1001111";--  -11
			when "011110110"=>x3<="1111110";x2<="0000001";x1<="1001111";x0<="0000001";--  -10
			when "011110111"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0001000";--  -9
			when "011111000"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0000000";--  -8
			when "011111001"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0001111";-- -7
			when "011111010"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0100000";-- -6
			when "011111011"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0100100";-- -5
			when "011111100"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="1001100";-- -4
			when "011111101"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0000110";-- -3
			when "011111110"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="0010010";-- -2
			when "011111111"=>x3<="1111110";x2<="0000001";x1<="0000001";x0<="1001111";-- -1	
			when others=>x3<="1001000";x2<="1001000";x1<="1001000";x0<="1001000"; -- H,codul de eroare 
		end case;																			 

		end process;
end f1;