library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
entity s is
end ;
architecture f of s is	 
 signal numar1:std_logic_vector(3 downto 0):=x"0";
begin

end ;